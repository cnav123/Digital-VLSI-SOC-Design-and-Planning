magic
tech sky130A
timestamp 1598787264
<< metal1 >>
rect 0 90 45 105
rect 30 0 45 90
<< properties >>
string FIXED_BBOX 0 -30 60 105
<< end >>
